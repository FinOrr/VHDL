library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity Channel_B is
    generic (
        LFSR_Seed    :  std_logic_vector(32 downto 1) := x"3CA52DF7"    -- Generic seed to intialise the PRNG
    );
    port (
        -- Inputs
        Clk          :  in  std_logic;                                  -- System clock
        Clock_En     :  in  std_logic;                                  -- Clock enable signal
        Reset        :  in  std_logic;                                  -- Global reset signal
        Error_Select :  in  std_logic_vector(1 downto 0);               -- 2 bit input to control the error to be introduced
        I_RX         :  in  std_logic_vector(7 downto 0);               -- Input of I channel
        Q_RX         :  in  std_logic_vector(7 downto 0);               -- Input of the Q channel
        
        -- Outputs
        I_TX         :  out std_logic_vector(7 downto 0);               -- I channel output, with random error
        Q_TX         :  out std_logic_vector(7 downto 0)                -- Q channel output, with random error
    );
end Channel_B;

architecture Behavioral of Channel_B is

    signal Error_Raw    : std_logic_vector(7 downto 0);                 -- Random error generated by taking values from LFSR
    signal Error_16     : std_logic_vector(7 downto 0);                 -- Random error, clamped to only give values between +- 16
    signal Error_32     : std_logic_vector(7 downto 0);                 -- Random error that only gives values between +- 32
    signal Error_64     : std_logic_vector(7 downto 0);                 -- Random error, clamped to only give values between +- 64
    signal LFSR         : std_logic_vector(32 downto 1) := LFSR_Seed;   -- Seed the LFSR
    signal XNOR_Bit     : std_logic := '0';
    
begin

    ----------------------------------------------------------------------------------
    --                      Generating the error signal                             --
    ----------------------------------------------------------------------------------
    -- Bit Index:   7       6      5       4      3       2       1       0         --
    -- Bit value:   +-      64     32      16     8       4       2       1         --
    --      NOTE: IF sign bit AND bit 6 = 0,              error value is < +64      --
    --            IF sign bit AND bit 6 AND 5 = 0,        error value is < +32      --
    --            IF sign bit AND bit 6 AND 5 AND 4  = 0, error value is < +16      --
    --                                                                              --
    --      NOTE: IF SIGN BIT = 1 (i.e the error is negative) then bits             --
    --            6, 5, 4 will need to be set to 1 instead of 0                     --
    ----------------------------------------------------------------------------------
    
    ---- Error introduction process 
    Error_Addition: process(Clk)
    begin
        if (rising_edge(Clk)) then            
            if (Clock_En = '1') then
        
            Error_Raw(7 downto 0) <= LFSR(32 downto 25);                 -- Values for the Error signal are pulled from the LFSR
            
            -- Bit mask error signals --
            if (Error_Raw(7) = '1') then                                 -- Check if the random error is a negative number
                Error_16(7 downto 0) <= "1111" & Error_Raw(3 downto 0);  -- Mask bits 4,5,6 with '1' so Error_16 is within the acceptable range when negative
                Error_32(7 downto 0) <= "111"  & Error_Raw(4 downto 0);  -- Mask bits 5 and 6 with '1' so Error_32 gives a maximum negative value of -32
                Error_64(7 downto 0) <= "11"   & Error_Raw(5 downto 0);  -- Mask bit 6 with a '1', so the most negative value of Error_64 is -64                    
            else
                Error_16(7 downto 0) <= "0000" & Error_Raw(3 downto 0);  -- Mask bits 4,5,6 with '0' so Error_16 is within the acceptable range when positive
                Error_32(7 downto 0) <= "000"  & Error_Raw(4 downto 0);  -- Mask bits 5 and 6 with '0' so Error_32 gives a maximum value of +31
                Error_64(7 downto 0) <= "00"   & Error_Raw(5 downto 0);  -- Mask bit 6 with a '0', so the greatest value of Error_64 is +63
            end if; -- end polarity check
                
            -- Case statement generates the output of the channel block depending on the error select input
            case Error_Select is
            
                when "00" =>        -- No Error
                    I_TX <= I_RX;
                    Q_TX <= Q_RX;
                
                when "01" =>        -- (+- 16 error)                        
                    I_TX <= std_logic_vector(unsigned(I_RX) + unsigned(Error_16));
                    Q_TX <= std_logic_vector(unsigned(I_RX) + unsigned(Error_16));
                
                when "10" =>        -- (+- 32 error)
                    I_TX <= std_logic_vector(unsigned(I_RX) + unsigned(Error_32));
                    Q_TX <= std_logic_vector(unsigned(I_RX) + unsigned(Error_32));
                    
                when "11" =>        -- (+- 64 error)
                    I_TX <= std_logic_vector(unsigned(I_RX) + unsigned(Error_64));
                    Q_TX <= std_logic_vector(unsigned(I_RX) + unsigned(Error_64));
                                            
                when others =>      -- others statement to catch errors
                    I_TX <= (others => 'Z');
                    Q_TX <= (others => 'Z');
                    
                end case; -- end error select check case
            end if; -- End clock enable check
        end if; -- end rising edge check 
    end process; -- end Error_Convolution process
    
    
    ---- Pseudo random number generator using a linear feedback shift register -----
    PRN_Generator: process(Clk)
    begin   
        if (rising_edge(Clk)) then                                              -- Sync on system clock
            if (Reset = '1') then                                               -- Check for synchronous reset
                LFSR <= LFSR_Seed;                                              -- If reset is true, reset LFSR to initial seed
            elsif (Clock_En = '1') then                                         -- Sync number generation to clock enable
                XNOR_Bit <= LFSR(32) xnor LFSR(22) xnor LFSR(2) xnor LFSR(1);   -- New bit to be shifted into LFSR is generated by XNOR'ing bits
                LFSR     <= LFSR(31 downto 1) & XNOR_Bit;                       -- Shift new bit into the LFSR
            end if;
        end if;
    end process;

end Behavioral;