library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package TYPES is

    type t_Waveform is array(7 downto 0) of std_logic_vector(7 downto 0);

end package;